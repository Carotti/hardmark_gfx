package vector;

    typedef struct packed {
        fixed_point::fixed_point_t x;
        fixed_point::fixed_point_t y;
        fixed_point::fixed_point_t z;
    } vector_t;

endpackage