package graphics;

    typedef struct packed {
        vector::vector_t intersection_point;
        logic intersects;
    } intersection_t;

endpackage