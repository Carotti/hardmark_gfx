package fixed_point;

    typedef struct packed {
        logic [18:0] i;
        logic [12:0] f; 
    } fixed_point_t;

endpackage